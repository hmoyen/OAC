module riscv_fd (
    input clock,
    input reset
);

    
endmodule