module riscv_uc (
    input clock,
    input reset
);

    
endmodule