module moduleName (
    input clock,
    input reset,
    input start,
    output done
);
    
riscv_uc UC (

);

riscv_fd FD (

);

endmodule